`include "../../sys_defs.vh"
module icache(
    input   clock,
    input   reset,
    input   [3:0] Imem2proc_response1,
    input   [3:0] Imem2proc_response ,
    input  [63:0] Imem2proc_data1,
    input  [63:0] Imem2proc_data,
    input   [3:0] Imem2proc_tag1,
    input   [3:0] Imem2proc_tag,

    input  [63:0] proc2Icache_addr1,
    input  [63:0] proc2Icache_addr,
    input  [63:0] cachemem_data1,
    input  [63:0] cachemem_data,
    input   cachemem_valid1,
    input   cachemem_valid,

    output logic  [1:0] proc2Imem_command1,
    output logic  [1:0] proc2Imem_command ,
    output logic [63:0] proc2Imem_addr1,
    output logic [63:0] proc2Imem_addr,

    output logic [63:0] Icache_data_out1, // value is memory[proc2Icache_addr]
    output logic [63:0] Icache_data_out, // value is memory[proc2Icache_addr]
    output logic  Icache_valid_out1,      // when this is high
    output logic  Icache_valid_out,      // when this is high

    output logic  [(`NUM_SET_BITS - 1):0] current_index1,
    output logic  [(`NUM_SET_BITS - 1):0] current_index,
    output logic  [(`NUM_TAG_BITS - 1):0] current_tag1,
    output logic  [(`NUM_TAG_BITS - 1):0] current_tag,
    output logic  [(`NUM_SET_BITS - 1):0] last_index1,
    output logic  [(`NUM_SET_BITS - 1):0] last_index,
    output logic  [(`NUM_TAG_BITS - 1):0] last_tag1,
    output logic  [(`NUM_TAG_BITS - 1):0] last_tag,
    output logic  data_write_enable1,
    output logic  data_write_enable
  
  );

  logic [3:0] current_mem_tag1;
  logic [3:0] current_mem_tag;

  logic miss_outstanding1;
  logic miss_outstanding;

  assign {current_tag1, current_index1} = proc2Icache_addr1[31:3];
  assign {current_tag , current_index } = proc2Icache_addr [31:3];

  wire changed_addr1 = (current_index1 != last_index1) || (current_tag1 != last_tag1);
  wire changed_addr  = (current_index  != last_index ) || (current_tag  != last_tag );

  wire send_request1 = miss_outstanding1 && !changed_addr1;
  wire send_request  = miss_outstanding  && !changed_addr ;

  assign Icache_data_out1 = cachemem_data1;
  assign Icache_data_out  = cachemem_data ;

  assign Icache_valid_out1 = cachemem_valid1; 
  assign Icache_valid_out  = cachemem_valid ; 

  assign proc2Imem_addr1 = {proc2Icache_addr1[63:3],3'b0};
  assign proc2Imem_addr  = {proc2Icache_addr [63:3],3'b0};
  assign proc2Imem_command1 = (miss_outstanding1 && !changed_addr1) ?  BUS_LOAD :
                                                                    BUS_NONE;
  assign proc2Imem_command  = (miss_outstanding  && !changed_addr ) ?  BUS_LOAD :
                                                                    BUS_NONE;                                                                  

 // assign data_write_enable =  (current_mem_tag == Imem2proc_tag) &&
                           //   (current_mem_tag != 0);
  assign data_write_enable1 = (Imem2proc_response1 == Imem2proc_tag1) && (Imem2proc_response1 != 0);
  assign data_write_enable  = (Imem2proc_response  == Imem2proc_tag ) && (Imem2proc_response  != 0);

  wire update_mem_tag1 = changed_addr1 || miss_outstanding1 || data_write_enable1;
  wire update_mem_tag  = changed_addr  || miss_outstanding  || data_write_enable ;

  wire unanswered_miss1 = changed_addr1 ? !Icache_valid_out1 :
                                        miss_outstanding1 && (Imem2proc_response1 == 0);
  wire unanswered_miss  = changed_addr  ? !Icache_valid_out  :
                                        miss_outstanding  && (Imem2proc_response  == 0);                                      

  // synopsys sync_set_reset "reset"
  always_ff @(posedge clock) begin
    if(reset) begin
      last_index1       <= `SD -1;   // These are -1 to get ball rolling when
      last_index        <= `SD -1;   // These are -1 to get ball rolling when
      last_tag1         <= `SD -1;   // reset goes low because addr "changes"
      last_tag          <= `SD -1;   // reset goes low because addr "changes"
      current_mem_tag1  <= `SD 0;
      current_mem_tag   <= `SD 0;              
      miss_outstanding1 <= `SD 0;
      miss_outstanding  <= `SD 0;
    end else begin
      last_index1       <= `SD current_index1;
      last_index        <= `SD current_index ;
      last_tag1         <= `SD current_tag1;
      last_tag          <= `SD current_tag ;
      miss_outstanding1 <= `SD unanswered_miss1;
      miss_outstanding  <= `SD unanswered_miss ;
      
      if(update_mem_tag1)
        current_mem_tag1 <= `SD Imem2proc_response1;
      if(update_mem_tag )
        current_mem_tag  <= `SD Imem2proc_response ;
    end
  end

endmodule


`include "../../sys_defs.vh"
`define DEBUG
`define DELAY #2
`define CLOCK_PERIOD #10
`define NUM_RAND_ITER 500

module testbench;

	initial
	begin
		$finish;
	end


endmodule

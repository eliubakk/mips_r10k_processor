module Map_Table(
	input	clock,
	input 	reset,
	input	enable,
	
);
endmodule // Map_Table